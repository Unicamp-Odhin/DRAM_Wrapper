module Wrapper #(
    parameter SYS_CLK_FREQ = 100_000_000
) (
    input  logic sys_clk,
    input  logic rst_n,
);
    
endmodule
